// asm file name: jalr.o
module instr_rom(
    input  logic clk, rst_n,
    input  logic [13:0] i_addr,
    output logic [31:0] o_data
);
    localparam  INSTR_CNT = 12'd61;
    
    wire [0:INSTR_CNT-1] [31:0] instr_rom_cell = {
        32'h00200193,    //0x00000000
        32'h00000293,    //0x00000004
        32'h00000317,    //0x00000008
        32'h01030313,    //0x0000000c
        32'h000302e7,    //0x00000010
        32'h0c00006f,    //0x00000014
        32'h00000317,    //0x00000018
        32'hffc30313,    //0x0000001c
        32'h0a629a63,    //0x00000020
        32'h00400193,    //0x00000024
        32'h00000213,    //0x00000028 
        32'h00000317,    //0x0000002c
        32'h01030313,    //0x00000030
        32'h000309e7,    //0x00000034
        32'h08301e63,    //0x00000038
        32'h00120213,    //0x0000003c
        32'h00200293,    //0x00000040
        32'hfe5214e3,    //0x00000044
        32'h00500193,    //0x00000048
        32'h00000213,    //0x0000004c
        32'h00000317,    //0x00000050
        32'h01430313,    //0x00000054
        32'h00000013,    //0x00000058
        32'h000309e7,    //0x0000005c
        32'h06301a63,    //0x00000060
        32'h00120213,    //0x00000064
        32'h00200293,    //0x00000068
        32'hfe5212e3,    //0x0000006c
        32'h00600193,    //0x00000070
        32'h00000213,    //0x00000074
        32'h00000317,    //0x00000078
        32'h01830313,    //0x0000007c
        32'h00000013,    //0x00000080
        32'h00000013,    //0x00000084
        32'h000309e7,    //0x00000088
        32'h04301463,    //0x0000008c
        32'h00120213,    //0x00000090
        32'h00200293,    //0x00000094
        32'hfe5210e3,    //0x00000098
        32'h00100293,    //0x0000009c
        32'h00000317,    //0x000000a0
        32'h01c30313,    //0x000000a4
        32'hffc30067,    //0x000000a8
        32'h00128293,    //0x000000ac
        32'h00128293,    //0x000000b0
        32'h00128293,    //0x000000b4
        32'h00128293,    //0x000000b8
        32'h00128293,    //0x000000bc
        32'h00128293,    //0x000000c0
        32'h00400e93,    //0x000000c4
        32'h00700193,    //0x000000c8
        32'h01d29463,    //0x000000cc
        32'h00301863,    //0x000000d0
        32'h00100793,    //0x000000d4
        32'h00000213,    //0x000000d8
        32'h00320233,    //0x000000dc
        32'h00100193,    //0x000000e0
        32'h40f181b3,    //0x000000e4
        32'hc0001073,    //0x000000e8
        32'h00000000,    //0x000000ec
        32'h00000000    //0x000000f0
    };
    
    logic [11:0] instr_index;
    logic [31:0] data;
    
    assign instr_index = i_addr[13:2];
    assign data = (instr_index>=INSTR_CNT) ? 0 : instr_rom_cell[instr_index];
    
    always @ (posedge clk or negedge rst_n)
        if(~rst_n)
            o_data <= 0;
        else
            o_data <= data;

endmodule
