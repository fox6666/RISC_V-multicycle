// asm file name: add.o
module instr_rom(
    input  logic clk, rst_n,
    input  logic [13:0] i_addr,
    output logic [31:0] o_data
);
    localparam  INSTR_CNT = 12'd321;
    
    wire [0:INSTR_CNT-1] [31:0] instr_rom_cell = {
        32'h00000093,    //0x00000000
        32'h00000113,    //0x00000004
        32'h00208f33,    //0x00000008
        32'h00000e93,    //0x0000000c
        32'h00200193,    //0x00000010
        32'h4ddf1663,    //0x00000014
        32'h00100093,    //0x00000018
        32'h00100113,    //0x0000001c
        32'h00208f33,    //0x00000020
        32'h00200e93,    //0x00000024
        32'h00300193,    //0x00000028
        32'h4bdf1a63,    //0x0000002c
        32'h00300093,    //0x00000030
        32'h00700113,    //0x00000034
        32'h00208f33,    //0x00000038
        32'h00a00e93,    //0x0000003c
        32'h00400193,    //0x00000040
        32'h49df1e63,    //0x00000044
        32'h00000093,    //0x00000048
        32'hffff8137,    //0x0000004c
        32'h00208f33,    //0x00000050
        32'hffff8eb7,    //0x00000054
        32'h00500193,    //0x00000058
        32'h49df1263,    //0x0000005c
        32'h800000b7,    //0x00000060
        32'h00000113,    //0x00000064
        32'h00208f33,    //0x00000068
        32'h80000eb7,    //0x0000006c
        32'h00600193,    //0x00000070
        32'h47df1663,    //0x00000074
        32'h800000b7,    //0x00000078
        32'hffff8137,    //0x0000007c
        32'h00208f33,    //0x00000080
        32'h7fff8eb7,    //0x00000084
        32'h00700193,    //0x00000088
        32'h45df1a63,    //0x0000008c
        32'h00000093,    //0x00000090
        32'h00008137,    //0x00000094
        32'hfff10113,    //0x00000098
        32'h00208f33,    //0x0000009c
        32'h00008eb7,    //0x000000a0
        32'hfffe8e93,    //0x000000a4
        32'h00800193,    //0x000000a8
        32'h43df1a63,    //0x000000ac
        32'h800000b7,    //0x000000b0
        32'hfff08093,    //0x000000b4
        32'h00000113,    //0x000000b8
        32'h00208f33,    //0x000000bc
        32'h80000eb7,    //0x000000c0
        32'hfffe8e93,    //0x000000c4
        32'h00900193,    //0x000000c8
        32'h41df1a63,    //0x000000cc
        32'h800000b7,    //0x000000d0
        32'hfff08093,    //0x000000d4
        32'h00008137,    //0x000000d8
        32'hfff10113,    //0x000000dc
        32'h00208f33,    //0x000000e0
        32'h80008eb7,    //0x000000e4
        32'hffee8e93,    //0x000000e8
        32'h00a00193,    //0x000000ec
        32'h3fdf1863,    //0x000000f0
        32'h800000b7,    //0x000000f4
        32'h00008137,    //0x000000f8
        32'hfff10113,    //0x000000fc
        32'h00208f33,    //0x00000100
        32'h80008eb7,    //0x00000104
        32'hfffe8e93,    //0x00000108
        32'h00b00193,    //0x0000010c
        32'h3ddf1863,    //0x00000110
        32'h800000b7,    //0x00000114
        32'hfff08093,    //0x00000118
        32'hffff8137,    //0x0000011c
        32'h00208f33,    //0x00000120
        32'h7fff8eb7,    //0x00000124
        32'hfffe8e93,    //0x00000128
        32'h00c00193,    //0x0000012c
        32'h3bdf1863,    //0x00000130
        32'h00000093,    //0x00000134
        32'hfff00113,    //0x00000138
        32'h00208f33,    //0x0000013c
        32'hfff00e93,    //0x00000140
        32'h00d00193,    //0x00000144
        32'h39df1c63,    //0x00000148
        32'hfff00093,    //0x0000014c
        32'h00100113,    //0x00000150
        32'h00208f33,    //0x00000154
        32'h00000e93,    //0x00000158
        32'h00e00193,    //0x0000015c
        32'h39df1063,    //0x00000160
        32'hfff00093,    //0x00000164
        32'hfff00113,    //0x00000168
        32'h00208f33,    //0x0000016c
        32'hffe00e93,    //0x00000170
        32'h00f00193,    //0x00000174
        32'h37df1463,    //0x00000178
        32'h00100093,    //0x0000017c
        32'h80000137,    //0x00000180
        32'hfff10113,    //0x00000184
        32'h00208f33,    //0x00000188
        32'h80000eb7,    //0x0000018c
        32'h01000193,    //0x00000190
        32'h35df1663,    //0x00000194
        32'h00d00093,    //0x00000198
        32'h00b00113,    //0x0000019c
        32'h002080b3,    //0x000001a0
        32'h01800e93,    //0x000001a4
        32'h01100193,    //0x000001a8
        32'h33d09a63,    //0x000001ac
        32'h00e00093,    //0x000001b0
        32'h00b00113,    //0x000001b4
        32'h00208133,    //0x000001b8
        32'h01900e93,    //0x000001bc
        32'h01200193,    //0x000001c0
        32'h31d11e63,    //0x000001c4
        32'h00d00093,    //0x000001c8
        32'h001080b3,    //0x000001cc
        32'h01a00e93,    //0x000001d0
        32'h01300193,    //0x000001d4
        32'h31d09463,    //0x000001d8
        32'h00000213,    //0x000001dc
        32'h00d00093,    //0x000001e0
        32'h00b00113,    //0x000001e4
        32'h00208f33,    //0x000001e8
        32'h000f0313,    //0x000001ec
        32'h00120213,    //0x000001f0
        32'h00200293,    //0x000001f4
        32'hfe5214e3,    //0x000001f8
        32'h01800e93,    //0x000001fc
        32'h01400193,    //0x00000200
        32'h2dd31e63,    //0x00000204
        32'h00000213,    //0x00000208
        32'h00e00093,    //0x0000020c
        32'h00b00113,    //0x00000210
        32'h00208f33,    //0x00000214
        32'h00000013,    //0x00000218
        32'h000f0313,    //0x0000021c
        32'h00120213,    //0x00000220
        32'h00200293,    //0x00000224
        32'hfe5212e3,    //0x00000228
        32'h01900e93,    //0x0000022c
        32'h01500193,    //0x00000230
        32'h2bd31663,    //0x00000234
        32'h00000213,    //0x00000238
        32'h00f00093,    //0x0000023c
        32'h00b00113,    //0x00000240
        32'h00208f33,    //0x00000244
        32'h00000013,    //0x00000248
        32'h00000013,    //0x0000024c
        32'h000f0313,    //0x00000250
        32'h00120213,    //0x00000254
        32'h00200293,    //0x00000258
        32'hfe5210e3,    //0x0000025c
        32'h01a00e93,    //0x00000260
        32'h01600193,    //0x00000264
        32'h27d31c63,    //0x00000268
        32'h00000213,    //0x0000026c
        32'h00d00093,    //0x00000270
        32'h00b00113,    //0x00000274
        32'h00208f33,    //0x00000278
        32'h00120213,    //0x0000027c
        32'h00200293,    //0x00000280
        32'hfe5216e3,    //0x00000284
        32'h01800e93,    //0x00000288
        32'h01700193,    //0x0000028c
        32'h25df1863,    //0x00000290
        32'h00000213,    //0x00000294
        32'h00e00093,    //0x00000298
        32'h00b00113,    //0x0000029c
        32'h00000013,    //0x000002a0
        32'h00208f33,    //0x000002a4
        32'h00120213,    //0x000002a8
        32'h00200293,    //0x000002ac
        32'hfe5214e3,    //0x000002b0
        32'h01900e93,    //0x000002b4
        32'h01800193,    //0x000002b8
        32'h23df1263,    //0x000002bc
        32'h00000213,    //0x000002c0
        32'h00f00093,    //0x000002c4
        32'h00b00113,    //0x000002c8
        32'h00000013,    //0x000002cc
        32'h00000013,    //0x000002d0
        32'h00208f33,    //0x000002d4
        32'h00120213,    //0x000002d8
        32'h00200293,    //0x000002dc
        32'hfe5212e3,    //0x000002e0
        32'h01a00e93,    //0x000002e4
        32'h01900193,    //0x000002e8
        32'h1fdf1a63,    //0x000002ec
        32'h00000213,    //0x000002f0
        32'h00d00093,    //0x000002f4
        32'h00000013,    //0x000002f8
        32'h00b00113,    //0x000002fc
        32'h00208f33,    //0x00000300
        32'h00120213,    //0x00000304
        32'h00200293,    //0x00000308
        32'hfe5214e3,    //0x0000030c
        32'h01800e93,    //0x00000310
        32'h01a00193,    //0x00000314
        32'h1ddf1463,    //0x00000318
        32'h00000213,    //0x0000031c
        32'h00e00093,    //0x00000320
        32'h00000013,    //0x00000324
        32'h00b00113,    //0x00000328
        32'h00000013,    //0x0000032c
        32'h00208f33,    //0x00000330
        32'h00120213,    //0x00000334
        32'h00200293,    //0x00000338
        32'hfe5212e3,    //0x0000033c
        32'h01900e93,    //0x00000340
        32'h01b00193,    //0x00000344
        32'h19df1c63,    //0x00000348
        32'h00000213,    //0x0000034c
        32'h00f00093,    //0x00000350
        32'h00000013,    //0x00000354
        32'h00000013,    //0x00000358
        32'h00b00113,    //0x0000035c
        32'h00208f33,    //0x00000360
        32'h00120213,    //0x00000364
        32'h00200293,    //0x00000368
        32'hfe5212e3,    //0x0000036c
        32'h01a00e93,    //0x00000370
        32'h01c00193,    //0x00000374
        32'h17df1463,    //0x00000378
        32'h00000213,    //0x0000037c
        32'h00b00113,    //0x00000380
        32'h00d00093,    //0x00000384
        32'h00208f33,    //0x00000388
        32'h00120213,    //0x0000038c
        32'h00200293,    //0x00000390
        32'hfe5216e3,    //0x00000394
        32'h01800e93,    //0x00000398
        32'h01d00193,    //0x0000039c
        32'h15df1063,    //0x000003a0
        32'h00000213,    //0x000003a4
        32'h00b00113,    //0x000003a8
        32'h00e00093,    //0x000003ac
        32'h00000013,    //0x000003b0
        32'h00208f33,    //0x000003b4
        32'h00120213,    //0x000003b8
        32'h00200293,    //0x000003bc
        32'hfe5214e3,    //0x000003c0
        32'h01900e93,    //0x000003c4
        32'h01e00193,    //0x000003c8
        32'h11df1a63,    //0x000003cc
        32'h00000213,    //0x000003d0
        32'h00b00113,    //0x000003d4
        32'h00f00093,    //0x000003d8
        32'h00000013,    //0x000003dc
        32'h00000013,    //0x000003e0
        32'h00208f33,    //0x000003e4
        32'h00120213,    //0x000003e8
        32'h00200293,    //0x000003ec
        32'hfe5212e3,    //0x000003f0
        32'h01a00e93,    //0x000003f4
        32'h01f00193,    //0x000003f8
        32'h0fdf1263,    //0x000003fc
        32'h00000213,    //0x00000400
        32'h00b00113,    //0x00000404
        32'h00000013,    //0x00000408
        32'h00d00093,    //0x0000040c
        32'h00208f33,    //0x00000410
        32'h00120213,    //0x00000414
        32'h00200293,    //0x00000418
        32'hfe5214e3,    //0x0000041c
        32'h01800e93,    //0x00000420
        32'h02000193,    //0x00000424
        32'h0bdf1c63,    //0x00000428
        32'h00000213,    //0x0000042c
        32'h00b00113,    //0x00000430
        32'h00000013,    //0x00000434
        32'h00e00093,    //0x00000438
        32'h00000013,    //0x0000043c
        32'h00208f33,    //0x00000440
        32'h00120213,    //0x00000444
        32'h00200293,    //0x00000448
        32'hfe5212e3,    //0x0000044c
        32'h01900e93,    //0x00000450
        32'h02100193,    //0x00000454
        32'h09df1463,    //0x00000458
        32'h00000213,    //0x0000045c
        32'h00b00113,    //0x00000460
        32'h00000013,    //0x00000464
        32'h00000013,    //0x00000468
        32'h00f00093,    //0x0000046c
        32'h00208f33,    //0x00000470
        32'h00120213,    //0x00000474
        32'h00200293,    //0x00000478
        32'hfe5212e3,    //0x0000047c
        32'h01a00e93,    //0x00000480
        32'h02200193,    //0x00000484
        32'h05df1c63,    //0x00000488
        32'h00f00093,    //0x0000048c
        32'h00100133,    //0x00000490
        32'h00f00e93,    //0x00000494
        32'h02300193,    //0x00000498
        32'h05d11263,    //0x0000049c
        32'h02000093,    //0x000004a0
        32'h00008133,    //0x000004a4
        32'h02000e93,    //0x000004a8
        32'h02400193,    //0x000004ac
        32'h03d11863,    //0x000004b0
        32'h000000b3,    //0x000004b4
        32'h00000e93,    //0x000004b8
        32'h02500193,    //0x000004bc
        32'h03d09063,    //0x000004c0
        32'h01000093,    //0x000004c4
        32'h01e00113,    //0x000004c8
        32'h00208033,    //0x000004cc
        32'h00000e93,    //0x000004d0
        32'h02600193,    //0x000004d4
        32'h01d01463,    //0x000004d8
        32'h00301663,    //0x000004dc
        32'h00100793,    //0x000004e0
        32'h00320233,    //0x000004e4
        32'h00100193,    //0x000004e8
        32'h40f181b3,    //0x000004ec
        32'hc0001073,    //0x000004f0
        32'h00000000,    //0x000004f4
        32'h00000000,    //0x000004f8
        32'h00000000,    //0x000004fc
        32'h00000000    //0x00000500

    };
    
    logic [11:0] instr_index;
    logic [31:0] data;
    
    assign instr_index = i_addr[13:2];
    assign data = (instr_index>=INSTR_CNT) ? 0 : instr_rom_cell[instr_index];
    
    always @ (posedge clk or negedge rst_n)
        if(~rst_n)
            o_data <= 0;
        else
            o_data <= data;

endmodule
